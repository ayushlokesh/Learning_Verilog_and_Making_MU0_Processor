// Verilog HDL for "COMP12111_lib", "display_decoder" "functional"
//
// COMP12111 Exercise 2 - Combinatorial Design
//
// Version 2022. P W Nutter
//
// This is the Verilog module for the display decoder
//
// The aim of this exercise is complete the combinatorial design
// for the alphanumeric display decoder. 
//
// DO NOT change the interface to this design or it may not be marked completely
// when submitted.
//
// Make sure you document your code and marks may be awarded/lost for the 
// quality of the comments given. Please document in the header the changes 
// made, when and by whom.
//
// Comments:

module display_decoder (input 		[3:0]  input_code,       // bcd input
			output reg 	[14:0] segment_pattern); // segment code output

// provide Verilog that described the required behaviour of the
// combinatorial design
// -----------------------------------------------------------------







endmodule  // end of module display_decoder

